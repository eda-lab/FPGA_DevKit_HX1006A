
module source_probe (
	source,
	probe);	

	output	[23:0]	source;
	input	[23:0]	probe;
endmodule
